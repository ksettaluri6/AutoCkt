Top level OpenLoop

.include "/tools/projects/ISG/isg_chips/projects/kourosh_DeepCkt/bag_workspace_GF14LPP/bag_deep_ckt/eval_engines/NGspice/ngspice_inputs/spice_models/45nm_bulk.txt"
.include "/tools/projects/ISG/isg_chips/projects/kourosh_DeepCkt/bag_workspace_GF14LPP/bag_deep_ckt/eval_engines/NGspice/ngspice_inputs/netlist/Nested_Gboosting/no_gb/ota.subckt"

Xota VDD 0 inp inn outp outn cm_ref i_ref OTA m_in=m_in m_tail=m_tail m_cas=m_cas m_csp=m_csp m_bias_ref_n=m_bias_ref_n m_bias_ref_p=m_bias_ref_p m_biasn_local_n=m_biasn_local_n m_biasn_local_p=m_biasn_local_p m_biasp_local_n=m_biasp_local_n m_biasp_local_p=m_biasp_local_p m_cmfb_tail=m_cmfb_tail m_cmfb_amp=m_cmfb_amp m_cmfb_load=m_cmfb_load
CL outp outn cload

* testbench specification
vVDD VDD 0 1.2
ibias VDD i_ref ibias

vin in 0 dc=0 ac=1.0
ein1 inp incm in 0 0.5
ein2 inn incm in 0 -0.5
vcm incm 0 dc=vicm
vcm_ref cm_ref 0 dc=vocm

* parameters
.param ibias=20u
.param vicm=0.9
.param vocm=0.6
.param cload=1p

* amp parameters
.param m_in=50 m_tail=10 m_cas=25 m_csp=50
* reference bias parameters
.param m_bias_ref_n=10 m_bias_ref_p=10
* loacl nmos bias parameters
.param m_biasn_local_n=10 m_biasn_local_p=10
* loacl pmos bias parameters
.param m_biasp_local_n=10 m_biasp_local_p=10
* cmfb parameters
.param m_cmfb_tail=10 m_cmfb_amp=10 m_cmfb_load=10


.ac dec 10 1 10G

.control
run
set units=degrees
set wr_vecnames
option numdgt=7
wrdata ac.csv v(outp)-v(outn)
op
wrdata dc.csv v(outp) v(outn) i(vVDD)
.endc

.end