** Generated for: hspiceD
** Generated on: Jan 24 07:27:35 2019
** Design library name: gain_boost_templates
** Design cell name: ac_tb
** Design view name: schematic
.PARAM ibais=20u m_bias_glob_n=2 m_bias_glob_p=4 m_bias_localn_n=2
+	m_bias_localn_p=4 m_bias_localp_n=2 m_bias_localp_p=4 m_main_csp=60
+	m_main_in=10 m_main_tail=10 vicm=900m vocm=0.6

.OPTION ARTIST=0 PSF=2
.AC DEC 10 1.0 100e9

.OP voltage 1

.TEMP 25.0
.OPTION
+    ARTIST=2
+    INGOLD=2
+    PARHIER=LOCAL
+    PSF=2
.LIB "/tools/gftech14/GF_PDK/14LPP-XL_V1.3.1.0/Models/HSPICE/models/LN14LPP_Hspice.lib" TT

** Library name: gain_boost_templates
** Cell name: core_n
** View name: schematic
.subckt core_n vdd vss cs_n cs_p gb_bot_inn gb_bot_inp gb_bot_outn gb_bot_outp gb_top_inn gb_top_inp gb_top_outn gb_top_outp in_minus in_plus o_minus o_plus tail_b tail_t
xmcs_n_l gb_bot_inn cs_n vss vss nfet m=1 l=14e-9 nfin=2 nf='(m_main_tail/2)*1' par=1 par_nf='1*((m_main_tail/2)*1)' asej='1.188e-15+(2*int((m_main_tail/2)/2))*594e-18' adej='(2*(1+int((m_main_tail/2-1)/2)))*594e-18' psej='227e-9+(((2*int((m_main_tail/2)/2))*1)*2)*54e-9' pdej='(((2*(1+int((m_main_tail/2-1)/2)))*1)*2)*54e-9' pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=38.988e-6 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xmcs_n_r gb_bot_inp cs_n vss vss nfet m=1 l=14e-9 nfin=2 nf='(m_main_tail/2)*1' par=1 par_nf='1*((m_main_tail/2)*1)' asej='1.188e-15+(2*int((m_main_tail/2)/2))*594e-18' adej='(2*(1+int((m_main_tail/2-1)/2)))*594e-18' psej='227e-9+(((2*int((m_main_tail/2)/2))*1)*2)*54e-9' pdej='(((2*(1+int((m_main_tail/2-1)/2)))*1)*2)*54e-9' pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=38.988e-6 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xmcas_n_l o_minus gb_bot_outp gb_bot_inn vss nfet m=1 l=14e-9 nfin=2 nf='(m_main_tail/2)*1' par=1 par_nf='1*((m_main_tail/2)*1)' asej='1.188e-15+(2*int((m_main_tail/2)/2))*594e-18' adej='(2*(1+int((m_main_tail/2-1)/2)))*594e-18' psej='227e-9+(((2*int((m_main_tail/2)/2))*1)*2)*54e-9' pdej='(((2*(1+int((m_main_tail/2-1)/2)))*1)*2)*54e-9' pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=38.988e-6 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xmcas_n_r o_plus gb_bot_outn gb_bot_inp vss nfet m=1 l=14e-9 nfin=2 nf='(m_main_tail/2)*1' par=1 par_nf='1*((m_main_tail/2)*1)' asej='1.188e-15+(2*int((m_main_tail/2)/2))*594e-18' adej='(2*(1+int((m_main_tail/2-1)/2)))*594e-18' psej='227e-9+(((2*int((m_main_tail/2)/2))*1)*2)*54e-9' pdej='(((2*(1+int((m_main_tail/2-1)/2)))*1)*2)*54e-9' pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=38.988e-6 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xmtail_bot net7 tail_b vss vss nfet m=1 l=14e-9 nfin=2 nf='m_main_tail*1' par=1 par_nf='1*(m_main_tail*1)' asej='1.188e-15+(2*int(m_main_tail/2))*594e-18' adej='(2*(1+int((m_main_tail-1)/2)))*594e-18' psej='227e-9+(((2*int(m_main_tail/2))*1)*2)*54e-9' pdej='(((2*(1+int((m_main_tail-1)/2)))*1)*2)*54e-9' pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=38.988e-6 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xmtail_top net1 tail_t net7 vss nfet m=1 l=14e-9 nfin=2 nf='m_main_tail*1' par=1 par_nf='1*(m_main_tail*1)' asej='1.188e-15+(2*int(m_main_tail/2))*594e-18' adej='(2*(1+int((m_main_tail-1)/2)))*594e-18' psej='227e-9+(((2*int(m_main_tail/2))*1)*2)*54e-9' pdej='(((2*(1+int((m_main_tail-1)/2)))*1)*2)*54e-9' pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=38.988e-6 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xmin_plus gb_top_inn in_plus net1 vss nfet m=1 l=14e-9 nfin=2 nf='m_main_in*1' par=1 par_nf='1*(m_main_in*1)' asej='1.188e-15+(2*int(m_main_in/2))*594e-18' adej='(2*(1+int((m_main_in-1)/2)))*594e-18' psej='227e-9+(((2*int(m_main_in/2))*1)*2)*54e-9' pdej='(((2*(1+int((m_main_in-1)/2)))*1)*2)*54e-9' pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=38.988e-6 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xmin_minus gb_top_inp in_minus net1 vss nfet m=1 l=14e-9 nfin=2 nf='m_main_in*1' par=1 par_nf='1*(m_main_in*1)' asej='1.188e-15+(2*int(m_main_in/2))*594e-18' adej='(2*(1+int((m_main_in-1)/2)))*594e-18' psej='227e-9+(((2*int(m_main_in/2))*1)*2)*54e-9' pdej='(((2*(1+int((m_main_in-1)/2)))*1)*2)*54e-9' pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=38.988e-6 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xmcas_p_l o_minus gb_top_outp gb_top_inn vdd pfet m=1 l=14e-9 nfin=2 nf='(m_main_csp/2)*1' par=1 par_nf='1*((m_main_csp/2)*1)' asej='1.188e-15+(2*int((m_main_csp/2)/2))*594e-18' adej='(2*(1+int((m_main_csp/2-1)/2)))*594e-18' psej='227e-9+(((2*int((m_main_csp/2)/2))*1)*2)*54e-9' pdej='(((2*(1+int((m_main_csp/2-1)/2)))*1)*2)*54e-9' pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=38.988e-6 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xmcs_p_l gb_top_inn cs_p vdd vdd pfet m=1 l=14e-9 nfin=2 nf='m_main_csp*1' par=1 par_nf='1*(m_main_csp*1)' asej='1.188e-15+(2*int(m_main_csp/2))*594e-18' adej='(2*(1+int((m_main_csp-1)/2)))*594e-18' psej='227e-9+(((2*int(m_main_csp/2))*1)*2)*54e-9' pdej='(((2*(1+int((m_main_csp-1)/2)))*1)*2)*54e-9' pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=38.988e-6 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xmcs_p_r gb_top_inp cs_p vdd vdd pfet m=1 l=14e-9 nfin=2 nf='m_main_csp*1' par=1 par_nf='1*(m_main_csp*1)' asej='1.188e-15+(2*int(m_main_csp/2))*594e-18' adej='(2*(1+int((m_main_csp-1)/2)))*594e-18' psej='227e-9+(((2*int(m_main_csp/2))*1)*2)*54e-9' pdej='(((2*(1+int((m_main_csp-1)/2)))*1)*2)*54e-9' pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=38.988e-6 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xmcas_p_r o_plus gb_top_outn gb_top_inp vdd pfet m=1 l=14e-9 nfin=2 nf='(m_main_csp/2)*1' par=1 par_nf='1*((m_main_csp/2)*1)' asej='1.188e-15+(2*int((m_main_csp/2)/2))*594e-18' adej='(2*(1+int((m_main_csp/2-1)/2)))*594e-18' psej='227e-9+(((2*int((m_main_csp/2)/2))*1)*2)*54e-9' pdej='(((2*(1+int((m_main_csp/2-1)/2)))*1)*2)*54e-9' pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=38.988e-6 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
.ends core_n
** End of subcircuit definition.

** Library name: gain_boost_templates
** Cell name: bias_global
** View name: schematic
.subckt bias_global vdd vss nb nt pb pt
xm5 pb pb pt vdd pfet m=1 l=14e-9 nfin=2 nf='m_bias_glob_p*1' par=1 par_nf='1*(m_bias_glob_p*1)' asej='1.188e-15+(2*int(m_bias_glob_p/2))*594e-18' adej='(2*(1+int((m_bias_glob_p-1)/2)))*594e-18' psej='227e-9+(((2*int(m_bias_glob_p/2))*1)*2)*54e-9' pdej='(((2*(1+int((m_bias_glob_p-1)/2)))*1)*2)*54e-9' pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=38.988e-6 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xm6 pt pt vdd vdd pfet m=1 l=14e-9 nfin=2 nf='m_bias_glob_p*1' par=1 par_nf='1*(m_bias_glob_p*1)' asej='1.188e-15+(2*int(m_bias_glob_p/2))*594e-18' adej='(2*(1+int((m_bias_glob_p-1)/2)))*594e-18' psej='227e-9+(((2*int(m_bias_glob_p/2))*1)*2)*54e-9' pdej='(((2*(1+int((m_bias_glob_p-1)/2)))*1)*2)*54e-9' pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=38.988e-6 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xm3 nb nb vss vss nfet m=1 l=14e-9 nfin=2 nf='m_bias_glob_n*1' par=1 par_nf='1*(m_bias_glob_n*1)' asej='1.188e-15+(2*int(m_bias_glob_n/2))*594e-18' adej='(2*(1+int((m_bias_glob_n-1)/2)))*594e-18' psej='227e-9+(((2*int(m_bias_glob_n/2))*1)*2)*54e-9' pdej='(((2*(1+int((m_bias_glob_n-1)/2)))*1)*2)*54e-9' pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=38.988e-6 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xm1 nt nt nb vss nfet m=1 l=14e-9 nfin=2 nf='m_bias_glob_n*1' par=1 par_nf='1*(m_bias_glob_n*1)' asej='1.188e-15+(2*int(m_bias_glob_n/2))*594e-18' adej='(2*(1+int((m_bias_glob_n-1)/2)))*594e-18' psej='227e-9+(((2*int(m_bias_glob_n/2))*1)*2)*54e-9' pdej='(((2*(1+int((m_bias_glob_n-1)/2)))*1)*2)*54e-9' pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=38.988e-6 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xm4 net14 nb vss vss nfet m=1 l=14e-9 nfin=2 nf='m_bias_glob_n*1' par=1 par_nf='1*(m_bias_glob_n*1)' asej='1.188e-15+(2*int(m_bias_glob_n/2))*594e-18' adej='(2*(1+int((m_bias_glob_n-1)/2)))*594e-18' psej='227e-9+(((2*int(m_bias_glob_n/2))*1)*2)*54e-9' pdej='(((2*(1+int((m_bias_glob_n-1)/2)))*1)*2)*54e-9' pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=38.988e-6 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xm2 pb nt net14 vss nfet m=1 l=14e-9 nfin=2 nf='m_bias_glob_n*1' par=1 par_nf='1*(m_bias_glob_n*1)' asej='1.188e-15+(2*int(m_bias_glob_n/2))*594e-18' adej='(2*(1+int((m_bias_glob_n-1)/2)))*594e-18' psej='227e-9+(((2*int(m_bias_glob_n/2))*1)*2)*54e-9' pdej='(((2*(1+int((m_bias_glob_n-1)/2)))*1)*2)*54e-9' pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=38.988e-6 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
.ends bias_global
** End of subcircuit definition.

** Library name: gain_boost_templates
** Cell name: bias_local_nmos
** View name: schematic
.subckt bias_local_nmos vdd vss nb nt pb pt
xm6 nb pb net15 vdd pfet m=1 l=14e-9 nfin=2 nf='m_bias_localn_p*1' par=1 par_nf='1*(m_bias_localn_p*1)' asej='1.188e-15+(2*int(m_bias_localn_p/2))*594e-18' adej='(2*(1+int((m_bias_localn_p-1)/2)))*594e-18' psej='227e-9+(((2*int(m_bias_localn_p/2))*1)*2)*54e-9' pdej='(((2*(1+int((m_bias_localn_p-1)/2)))*1)*2)*54e-9' pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=38.988e-6 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xm8 net15 pt vdd vdd pfet m=1 l=14e-9 nfin=2 nf='m_bias_localn_p*1' par=1 par_nf='1*(m_bias_localn_p*1)' asej='1.188e-15+(2*int(m_bias_localn_p/2))*594e-18' adej='(2*(1+int((m_bias_localn_p-1)/2)))*594e-18' psej='227e-9+(((2*int(m_bias_localn_p/2))*1)*2)*54e-9' pdej='(((2*(1+int((m_bias_localn_p-1)/2)))*1)*2)*54e-9' pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=38.988e-6 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xm5 nt pb net16 vdd pfet m=1 l=14e-9 nfin=2 nf='m_bias_localn_p*1' par=1 par_nf='1*(m_bias_localn_p*1)' asej='1.188e-15+(2*int(m_bias_localn_p/2))*594e-18' adej='(2*(1+int((m_bias_localn_p-1)/2)))*594e-18' psej='227e-9+(((2*int(m_bias_localn_p/2))*1)*2)*54e-9' pdej='(((2*(1+int((m_bias_localn_p-1)/2)))*1)*2)*54e-9' pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=38.988e-6 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xm7 net16 pt vdd vdd pfet m=1 l=14e-9 nfin=2 nf='m_bias_localn_p*1' par=1 par_nf='1*(m_bias_localn_p*1)' asej='1.188e-15+(2*int(m_bias_localn_p/2))*594e-18' adej='(2*(1+int((m_bias_localn_p-1)/2)))*594e-18' psej='227e-9+(((2*int(m_bias_localn_p/2))*1)*2)*54e-9' pdej='(((2*(1+int((m_bias_localn_p-1)/2)))*1)*2)*54e-9' pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=38.988e-6 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xm2 net13 nb vss vss nfet m=1 l=14e-9 nfin=2 nf='m_bias_localn_n*1' par=1 par_nf='1*(m_bias_localn_n*1)' asej='1.188e-15+(2*int(m_bias_localn_n/2))*594e-18' adej='(2*(1+int((m_bias_localn_n-1)/2)))*594e-18' psej='227e-9+(((2*int(m_bias_localn_n/2))*1)*2)*54e-9' pdej='(((2*(1+int((m_bias_localn_n-1)/2)))*1)*2)*54e-9' pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=38.988e-6 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xm4 nb nt net13 vss nfet m=1 l=14e-9 nfin=2 nf='m_bias_localn_n*1' par=1 par_nf='1*(m_bias_localn_n*1)' asej='1.188e-15+(2*int(m_bias_localn_n/2))*594e-18' adej='(2*(1+int((m_bias_localn_n-1)/2)))*594e-18' psej='227e-9+(((2*int(m_bias_localn_n/2))*1)*2)*54e-9' pdej='(((2*(1+int((m_bias_localn_n-1)/2)))*1)*2)*54e-9' pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=38.988e-6 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xm1 net14 nt vss vss nfet m=1 l=14e-9 nfin=2 nf='(m_bias_localn_n/2)*1' par=1 par_nf='1*((m_bias_localn_n/2)*1)' asej='1.188e-15+(2*int((m_bias_localn_n/2)/2))*594e-18' adej='(2*(1+int((m_bias_localn_n/2-1)/2)))*594e-18' psej='227e-9+(((2*int((m_bias_localn_n/2)/2))*1)*2)*54e-9' pdej='(((2*(1+int((m_bias_localn_n/2-1)/2)))*1)*2)*54e-9' pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=38.988e-6 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xm3 nt nt net14 vss nfet m=1 l=14e-9 nfin=2 nf='(m_bias_localn_n/2)*1' par=1 par_nf='1*((m_bias_localn_n/2)*1)' asej='1.188e-15+(2*int((m_bias_localn_n/2)/2))*594e-18' adej='(2*(1+int((m_bias_localn_n/2-1)/2)))*594e-18' psej='227e-9+(((2*int((m_bias_localn_n/2)/2))*1)*2)*54e-9' pdej='(((2*(1+int((m_bias_localn_n/2-1)/2)))*1)*2)*54e-9' pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=38.988e-6 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
.ends bias_local_nmos
** End of subcircuit definition.

** Library name: gain_boost_templates
** Cell name: bias_local_pmos
** View name: schematic
.subckt bias_local_pmos vdd vss nb nt pb pt
xm3 pb nt net15 vss nfet m=1 l=14e-9 nfin=2 nf='m_bias_localp_n*1' par=1 par_nf='1*(m_bias_localp_n*1)' asej='1.188e-15+(2*int(m_bias_localp_n/2))*594e-18' adej='(2*(1+int((m_bias_localp_n-1)/2)))*594e-18' psej='227e-9+(((2*int(m_bias_localp_n/2))*1)*2)*54e-9' pdej='(((2*(1+int((m_bias_localp_n-1)/2)))*1)*2)*54e-9' pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=38.988e-6 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xm1 net15 nb vss vss nfet m=1 l=14e-9 nfin=2 nf='m_bias_localp_n*1' par=1 par_nf='1*(m_bias_localp_n*1)' asej='1.188e-15+(2*int(m_bias_localp_n/2))*594e-18' adej='(2*(1+int((m_bias_localp_n-1)/2)))*594e-18' psej='227e-9+(((2*int(m_bias_localp_n/2))*1)*2)*54e-9' pdej='(((2*(1+int((m_bias_localp_n-1)/2)))*1)*2)*54e-9' pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=38.988e-6 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xm2 net16 nb vss vss nfet m=1 l=14e-9 nfin=2 nf='m_bias_localp_n*1' par=1 par_nf='1*(m_bias_localp_n*1)' asej='1.188e-15+(2*int(m_bias_localp_n/2))*594e-18' adej='(2*(1+int((m_bias_localp_n-1)/2)))*594e-18' psej='227e-9+(((2*int(m_bias_localp_n/2))*1)*2)*54e-9' pdej='(((2*(1+int((m_bias_localp_n-1)/2)))*1)*2)*54e-9' pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=38.988e-6 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xm4 pt nt net16 vss nfet m=1 l=14e-9 nfin=2 nf='m_bias_localp_n*1' par=1 par_nf='1*(m_bias_localp_n*1)' asej='1.188e-15+(2*int(m_bias_localp_n/2))*594e-18' adej='(2*(1+int((m_bias_localp_n-1)/2)))*594e-18' psej='227e-9+(((2*int(m_bias_localp_n/2))*1)*2)*54e-9' pdej='(((2*(1+int((m_bias_localp_n-1)/2)))*1)*2)*54e-9' pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=38.988e-6 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xm8 net13 pt vdd vdd pfet m=1 l=14e-9 nfin=2 nf='m_bias_localp_p*1' par=1 par_nf='1*(m_bias_localp_p*1)' asej='1.188e-15+(2*int(m_bias_localp_p/2))*594e-18' adej='(2*(1+int((m_bias_localp_p-1)/2)))*594e-18' psej='227e-9+(((2*int(m_bias_localp_p/2))*1)*2)*54e-9' pdej='(((2*(1+int((m_bias_localp_p-1)/2)))*1)*2)*54e-9' pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=38.988e-6 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xm6 pt pb net13 vdd pfet m=1 l=14e-9 nfin=2 nf='m_bias_localp_p*1' par=1 par_nf='1*(m_bias_localp_p*1)' asej='1.188e-15+(2*int(m_bias_localp_p/2))*594e-18' adej='(2*(1+int((m_bias_localp_p-1)/2)))*594e-18' psej='227e-9+(((2*int(m_bias_localp_p/2))*1)*2)*54e-9' pdej='(((2*(1+int((m_bias_localp_p-1)/2)))*1)*2)*54e-9' pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=38.988e-6 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xm7 net14 pb vdd vdd pfet m=1 l=14e-9 nfin=2 nf='(m_bias_localp_p/2)*1' par=1 par_nf='1*((m_bias_localp_p/2)*1)' asej='1.188e-15+(2*int((m_bias_localp_p/2)/2))*594e-18' adej='(2*(1+int((m_bias_localp_p/2-1)/2)))*594e-18' psej='227e-9+(((2*int((m_bias_localp_p/2)/2))*1)*2)*54e-9' pdej='(((2*(1+int((m_bias_localp_p/2-1)/2)))*1)*2)*54e-9' pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=38.988e-6 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xm5 pb pb net14 vdd pfet m=1 l=14e-9 nfin=2 nf='(m_bias_localp_p/2)*1' par=1 par_nf='1*((m_bias_localp_p/2)*1)' asej='1.188e-15+(2*int((m_bias_localp_p/2)/2))*594e-18' adej='(2*(1+int((m_bias_localp_p/2-1)/2)))*594e-18' psej='227e-9+(((2*int((m_bias_localp_p/2)/2))*1)*2)*54e-9' pdej='(((2*(1+int((m_bias_localp_p/2-1)/2)))*1)*2)*54e-9' pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=38.988e-6 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
.ends bias_local_pmos
** End of subcircuit definition.

** Library name: gain_boost_templates
** Cell name: core_p
** View name: schematic
.subckt core_p vdd vss cs_n cs_p gb_bot_inn gb_bot_inp gb_bot_outn gb_bot_outp gb_top_inn gb_top_inp gb_top_outn gb_top_outp in_minus in_plus o_minus o_plus tail_b tail_t
xmcas_n_l o_minus gb_bot_outp gb_bot_inn vss nfet m=1 l=14e-9 nfin=2 nf=1 par=1 par_nf=1 asej=1.188e-15 adej=1.188e-15 psej=238e-9 pdej=238e-9 pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=27e-9 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xmcas_n_r o_plus gb_bot_outn gb_bot_inp vss nfet m=1 l=14e-9 nfin=2 nf=1 par=1 par_nf=1 asej=1.188e-15 adej=1.188e-15 psej=238e-9 pdej=238e-9 pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=27e-9 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xmcs_n_l gb_bot_inn cs_n vss vss nfet m=1 l=14e-9 nfin=2 nf=1 par=1 par_nf=1 asej=1.188e-15 adej=1.188e-15 psej=238e-9 pdej=238e-9 pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=27e-9 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xmcs_n_r gb_bot_inp cs_n vss vss nfet m=1 l=14e-9 nfin=2 nf=1 par=1 par_nf=1 asej=1.188e-15 adej=1.188e-15 psej=238e-9 pdej=238e-9 pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=27e-9 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xmcs_p_l gb_top_inn cs_p vdd vdd pfet m=1 l=14e-9 nfin=2 nf=1 par=1 par_nf=1 asej=1.188e-15 adej=1.188e-15 psej=238e-9 pdej=238e-9 pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=27e-9 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xmcs_p_r gb_top_inp cs_p vdd vdd pfet m=1 l=14e-9 nfin=2 nf=1 par=1 par_nf=1 asej=1.188e-15 adej=1.188e-15 psej=238e-9 pdej=238e-9 pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=27e-9 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xmcas_p_l o_minus gb_top_outp gb_top_inn vdd pfet m=1 l=14e-9 nfin=2 nf=1 par=1 par_nf=1 asej=1.188e-15 adej=1.188e-15 psej=238e-9 pdej=238e-9 pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=27e-9 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xmcas_p_r o_plus gb_top_outn gb_top_inp vdd pfet m=1 l=14e-9 nfin=2 nf=1 par=1 par_nf=1 asej=1.188e-15 adej=1.188e-15 psej=238e-9 pdej=238e-9 pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=27e-9 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xmin_minus gb_bot_inp in_minus net7 vdd pfet m=1 l=14e-9 nfin=2 nf=1 par=1 par_nf=1 asej=1.188e-15 adej=1.188e-15 psej=238e-9 pdej=238e-9 pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=27e-9 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xmtail_top net16 tail_t vdd vdd pfet m=1 l=14e-9 nfin=2 nf=1 par=1 par_nf=1 asej=1.188e-15 adej=1.188e-15 psej=238e-9 pdej=238e-9 pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=27e-9 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xmtail_bot net7 tail_b net16 vdd pfet m=1 l=14e-9 nfin=2 nf=1 par=1 par_nf=1 asej=1.188e-15 adej=1.188e-15 psej=238e-9 pdej=238e-9 pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=27e-9 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
xmin_plus gb_bot_inn in_plus net7 vdd pfet m=1 l=14e-9 nfin=2 nf=1 par=1 par_nf=1 asej=1.188e-15 adej=1.188e-15 psej=238e-9 pdej=238e-9 pdevdops=1 pdevlgeos=1 pdevwgeos=1 psw_acv_sign=1 plnest=1 pldist=1 plorient=0 cpp=78e-9 fpitch=48e-9 xpos=-99 ypos=-99 ptwell=0 sca=0 scb=0 scc=0 pre_layout_local=-1 ngcon=1 p_vta=0 p_la=0 u0mult_fet=1 lle_sa=71e-9 lle_sb=71e-9 lle_rxrxa=78e-9 lle_rxrxb=78e-9 lle_rxrxn=192e-9 lle_rxrxs=192e-9 lle_pcrxn=65e-9 lle_pcrxs=65e-9 lle_nwa=2e-6 lle_nwb=2e-6 lle_nwn=192e-9 lle_nws=192e-9 lle_ctne=0 lle_ctnw=0 lle_ctse=0 lle_ctsw=0 lle_sctne=0 lle_sctnw=0 lle_sctse=0 lle_sctsw=0 lrsd=27e-9 dtemp=0 l_shape=0 l_shape_s=0 nsig_dop1=0 nsig_dop2=0 nsig_dibl=0 nsig_pc=0 nsig_rx=0 fc_index=0 fc_sigma=3
.ends core_p
** End of subcircuit definition.

** Library name: gain_boost_templates
** Cell name: folded_cascode_two_stage_gb
** View name: schematic
.subckt folded_cascode_two_stage_gb vdd vss i_ref in_minus in_plus o_minus o_plus vcm
xi31 vdd vss cs_n_b gb_bot_top_cmfb net023 net024 cs_n_t cs_n_t net025 net026 cs_p_b cs_p_b gb_bot_top_inn gb_bot_top_inp gb_bot_top_outn gb_bot_top_outp cs_n_b cs_n_t core_n
xi21 vdd vss cs_n_b gb_top_top_cmfb net014 net015 cs_n_t cs_n_t net013 net016 cs_p_b cs_p_b gb_top_top_inn gb_top_top_inp gb_top_top_outn gb_top_top_outp cs_n_b cs_n_t core_n
xgb1_top vdd vss cs_n_b gb_top_cmfb gb_top_bot_inn gb_top_bot_inp gb_top_bot_outn gb_top_bot_outp gb_top_top_inn gb_top_top_inp gb_top_top_outn gb_top_top_outp gb_top_inn gb_top_inp gb_top_outn gb_top_outp cs_n_b cs_n_t core_n
xcore_n vdd vss cs_n_b cmfb_minus gb_bot_inn gb_bot_inp gb_bot_outn gb_bot_outp gb_top_inn gb_top_inp gb_top_outn gb_top_outp in_minus in_plus o_minus o_plus cs_n_b cs_n_t core_n
xi0 vdd vss nb i_ref pb pt bias_global
xnmos_bias vdd vss cs_n_b cs_n_t pb pt bias_local_nmos
xpmos_bias vdd vss nb i_ref cs_p_b cs_p_t bias_local_pmos
e5 gb_bot_bot_cmfb vss VCVS gb_bot_bot_cm_out vcm 30
e4 gb_bot_top_cmfb vss VCVS gb_bot_top_cm_out vcm 30
e3 gb_top_bot_cmfb vss VCVS gb_top_bot_cm_out vcm 30
e2 gb_top_top_cmfb vss VCVS gb_top_top_cm_out vcm 30
e1 gb_bot_cmfb vss VCVS gb_bot_cm_out vcm 30
e0 gb_top_cmfb vss VCVS gb_top_cm_out vcm 30
evcmfb cmfb_minus vss VCVS cm_out vcm 30
r13 gb_bot_bot_outp gb_bot_bot_cm_out 1e12
r12 gb_bot_top_outn gb_bot_top_cm_out 1e12
r11 gb_bot_top_outp gb_bot_top_cm_out 1e12
r10 gb_bot_bot_outn gb_bot_bot_cm_out 1e12
r9 gb_top_bot_outp gb_top_bot_cm_out 1e12
r8 gb_top_bot_outn gb_top_bot_cm_out 1e12
r7 gb_top_top_outn gb_top_top_cm_out 1e12
r6 gb_top_top_outp gb_top_top_cm_out 1e12
r5 gb_bot_outp gb_bot_cm_out 1e12
r4 gb_bot_outn gb_bot_cm_out 1e12
r3 gb_top_outn gb_top_cm_out 1e12
r2 gb_top_outp gb_top_cm_out 1e12
r1 o_minus cm_out 1e12
r0 o_plus cm_out 1e12
c6 gb_bot_top_cm_out vss 1
c5 gb_bot_bot_cm_out vss 1
c4 gb_top_bot_cm_out vss 1
c3 gb_top_top_cm_out vss 1
c2 gb_bot_cm_out vss 1
c1 gb_top_cm_out vss 1
c0 cm_out vss 1
xi36 vdd vss gb_bot_bot_cmfb cs_p_t net029 net039 cs_n_t cs_n_t net030 net040 cs_p_b cs_p_b gb_bot_bot_inn gb_bot_bot_inp gb_bot_bot_outn gb_bot_bot_outp cs_p_b cs_p_t core_p
xi26 vdd vss gb_top_bot_cmfb cs_p_t net018 net027 cs_n_t cs_n_t net017 net028 cs_p_b cs_p_b gb_top_bot_inn gb_top_bot_inp gb_top_bot_outn gb_top_bot_outp cs_p_b cs_p_t core_p
xgb1_b vdd vss gb_bot_cmfb cs_p_t gb_bot_bot_inn gb_bot_bot_inp gb_bot_bot_outn gb_bot_bot_outp gb_bot_top_inn gb_bot_top_inp gb_bot_top_outn gb_bot_top_outp gb_bot_inn gb_bot_inp gb_bot_outn gb_bot_outp cs_p_b cs_p_t core_p
.ends folded_cascode_two_stage_gb
** End of subcircuit definition.

** Library name: gain_boost_templates
** Cell name: ac_tb
** View name: schematic
v11 in 0 DC=0 AC 1
v7 incm 0 DC=vicm
v1 vcm 0 DC=vocm
v0 vdd 0 DC=1.2
e3 in_plus incm VCVS in 0 -500e-3
e2 in_minus incm VCVS in 0 500e-3
i3 vdd i_ref DC=ibais
c0 o_plus o_minus 500e-15
xdut vdd 0 i_ref in_minus in_plus o_minus o_plus vcm folded_cascode_two_stage_gb
.END
